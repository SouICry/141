module CPU(
  input         start,
  input         CLK,
  output        halt);
  
  
endmodule